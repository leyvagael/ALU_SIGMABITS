LIBRARY IEEE;
USE ieee.std_logic_1164.all;

ENTITY FULL_ADDER IS
	PORT(
	A,B,Cin : IN STD_LOGIC;
	Co,S : OUT STD_LOGIC
	);
END FULL_ADDER;

ARCHITECTURE STRUCTURAL OF FULL_ADDER IS

COMPONENT HALF_ADDER
	PORT(
	A,B : IN STD_LOGIC;
	S,C : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL B0, B1, B2 : STD_LOGIC;

BEGIN
U0 : HALF_ADDER PORT MAP (A, B, B1, B0);
U1: HALF_ADDER PORT MAP (B1, Cin, S, B2);
Co <= B0 or B2;

END STRUCTURAL;